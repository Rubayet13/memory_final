`include "memory_packet.sv"
`include "memory_rtl.svp"
`include "memory_interface.sv"
`include "memory_driver.sv"
`include "memory_monitor.sv"
`include "memory_agent.sv"
`include "memory_scoreboard.sv"
`include "memory_env.sv"
`include "memory_test.sv"