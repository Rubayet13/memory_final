class packet;
	logic [7:0] data;
	logic [7:0] addr;


endclass  
